module memoryController
#(
	parameter S = 32,
	parameter V = 192,
	parameter SIZE_INS = 1000,
	parameter SIZE_ROM = 30000,
	parameter SIZE_RAM = 30000
)
(
);

endmodule