module mux_2to1_tb ();
	
	logic clk;
	logic [31:0] A, B, C, D, SAL1;
	logic [191:0] F, G, H, I, SAL2, SAL3, SAL4;
	logic sel;
	
	mux_2to1 #(32,32,32) mux_2to1_SSS (A, B, sel, SAL1);
	mux_2to1 #(32,192,192) mux_2to1_SVV (C, F, sel, SAL2);
	mux_2to1 #(192,32,192) mux_2to1_VSV (G, D, sel, SAL3);
	mux_2to1 #(192,192,192) mux_2to1_VVV (H, I, sel, SAL4);
	
	initial begin
		
		clk = 0; #2;
		
		// Mux 2 to 1, test 1:
		A = 32'b11110000111100001111000011110000; 
		B = 32'b11111111111111111111111111111111; 
		C = 32'b11111111111111111111111111111111;
		D = 32'b11111111111111111111111111111111;
		F = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		G = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		H = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		I = 192'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		sel = 1'b0; 
		#2;
		
		// Mux 2 to 1, test 2:
		A = 32'b11110000111100001111000011110000; 
		B = 32'b11111111111111111111111111111111; 
		C = 32'b11111111111111111111111111111111;
		D = 32'b11111111111111111111111111111111;
		F = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		G = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		H = 192'b100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001; 
		I = 192'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		sel = 1'b1; 
		#2;
		
	end
	
	always begin
		clk=!clk; #1;
	end
	
endmodule